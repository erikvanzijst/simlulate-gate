
* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create a pulse for A 
Va A VGND pulse(0 1.8 100p 10p 10p 100p 200p)

* setup the transient analysis
.tran 1p 3n 0

.control
run
set color0 = white
set color1 = black
plot A Y
.endc

.end
